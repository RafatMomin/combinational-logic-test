-- mux2t1_N.vhd (Structural)
library IEEE;
use IEEE.std_logic_1164.all;

entity mux2t1_N is
    generic(N : integer := 4); -- Default width set to 4
    port(
        i_S  : in std_logic;
        i_D0 : in std_logic_vector(N-1 downto 0);
        i_D1 : in std_logic_vector(N-1 downto 0);
        o_O  : out std_logic_vector(N-1 downto 0)
    );
end mux2t1_N;

architecture structural of mux2t1_N is

    -- Declare the mux2t1 component
    component mux2t1 is
        port(i_S    : in std_logic;
             i_D0   : in std_logic;
             i_D1   : in std_logic;
             o_O    : out std_logic);
    end component;

    -- Internal signals
    signal and_out0 : std_logic_vector(N-1 downto 0);
    signal and_out1 : std_logic_vector(N-1 downto 0);

begin
    -- Instantiate N-bit wide mux by instantiating 1-bit mux N times
    G_NBit_MUX: for i in 0 to N-1 generate
        MUXI: mux2t1
            port map(
                i_S    => i_S,
                i_D0   => i_D0(i),
                i_D1   => i_D1(i),
                o_O    => o_O(i)
            );
    end generate G_NBit_MUX;

end structural;