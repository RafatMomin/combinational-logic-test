library IEEE;
use IEEE.std_logic_1164.all;

entity tb_OnesComplementor is
    -- Testbench has no ports
end tb_OnesComplementor;

architecture behavior of tb_OnesComplementor is
    constant N : integer := 32;
    signal tb_i_A : std_logic_vector(N-1 downto 0);
    signal tb_o_F : std_logic_vector(N-1 downto 0);

    -- Instantiate the One's Complementor
begin
    uut: entity work.OnesComplementor
        generic map (N => N)
        port map (
            i_A => tb_i_A,
            o_F => tb_o_F
        );

    -- Process to apply test vectors and check results
    process
        -- Explicitly define expected output for each test case
        variable expected_all_zeros : std_logic_vector(N-1 downto 0) := (others => '1');
        variable expected_all_ones : std_logic_vector(N-1 downto 0) := (others => '0');
    begin
        -- Test vector 1: All zeros
        tb_i_A <= (others => '0');
        wait for 10 ns;
        assert tb_o_F = expected_all_zeros 
            --report "Test failed for all zeros input: Expected all ones, got " & std_logic_vector'image(tb_o_F)
            severity error;

        -- Test vector 2: All ones
        tb_i_A <= (others => '1');
        wait for 10 ns;
        assert tb_o_F = expected_all_ones 
           -- report "Test failed for all ones input: Expected all zeros, got " & std_logic_vector'image(tb_o_F)
            severity error;

        -- Test ends
        wait;
    end process;
end behavior;

